







    



    


                 


                 

                        





  





    

    



    

  







      





















                              ****** ********    ***********************                                             ****                ********************************












     





  *****************    
    
    
    
****            ****    ****                  

      







    






************                           
   
  
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    



  

          

                                       







      

      ****            
    
    
                                             

      

      

      

                              *******************************************************************                                                                                                                                                                                

                                                                                                
   ***************************************************************************                         **************************************************    ****                                                                                                                                                                                                                                                                                                                       						                                              														              																																																																																																																				                                               																															                                                                                                                                                                                                                                                                                                                                                                                                                                                                      																									      																																										                                                                                                                                                                                           													                                                          				                           	                																																																																																												         													                           																																																			                                                                                                                                                                                                                                                                                                                                                                                                        																					   										    												   				   						   																		   																																											                           															                       						                                                                       								    						       																														                                                                                                            																					    																								                                                                                            	                                                                                                                                                                                                                                    																																		         																																									 																																																					     																																																																																																																																																																										  									        													                                      			                                                                    						   								   						          																																										   													     																																																																																																					                                                                                                                                                             																																										        																																																															    			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           														                                                                                                                                                                             																																																																																				   						       			   																										       																																																																																																		   																																																                      			  																																																																																																																																								             									   									          																																																													                              																																																												 																																																																											                                             																																																																																																										     																					                                                         							 																								     																										                                       	                                                                                                                                                                                           																																       																																																																															               																																      				                            																																																																																																																	                     																	     																					                                                         				 							                                                                                                                       																																																													                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    .................           ..................                          .........................................                                                  ....                                      